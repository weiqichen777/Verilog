module fa(a, b, ci, sum, cout);
// input and output declaration
input  a, b, ci;
output sum, cout;

// wire and reg declaration


// module instance


endmodule

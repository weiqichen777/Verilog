// Serial Input BitStream Pattern Detector
module fsm_bspd(clk, reset, bit_in, det_out);
input clk, reset, bit_in;
output det_out;








endmodule

